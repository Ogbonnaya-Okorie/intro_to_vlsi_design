*** SPICE deck for cell r_divider_sim{sch} from library lab_1_dac
*** Created on Thu Sep 25, 2025 17:38:06
*** Last revised on Fri Sep 26, 2025 09:45:01
*** Written on Fri Sep 26, 2025 09:45:13 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT lab_1_dac__r_divider FROM CELL r_divider{sch}
.SUBCKT lab_1_dac__r_divider bot in out
Rresnwell@0 net@11 in 10k
Rresnwell@2 out bot 10k
Rresnwell@3 out net@11 10k
.ENDS lab_1_dac__r_divider

.global gnd

*** TOP LEVEL CELL: r_divider_sim{sch}
Xr_divide@0 gnd vin vout lab_1_dac__r_divider

* Spice Code nodes in cell cell 'r_divider_sim{sch}'
vin vin 0 DC 1
.op
.END
