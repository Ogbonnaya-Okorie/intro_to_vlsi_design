*** SPICE deck for cell dac_load_sim{sch} from library lab_1_dac
*** Created on Fri Sep 26, 2025 10:16:34
*** Last revised on Sun Sep 28, 2025 19:06:23
*** Written on Sun Sep 28, 2025 20:16:12 by Electric VLSI Design System, version 9.08
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT lab_1_dac__r_divider FROM CELL r_divider{sch}
.SUBCKT lab_1_dac__r_divider bot in out
Rresnwell@0 net@11 in 10k
Rresnwell@2 out bot 10k
Rresnwell@3 out net@11 10k
.ENDS lab_1_dac__r_divider

*** SUBCIRCUIT lab_1_dac__dac FROM CELL dac{sch}
.SUBCKT lab_1_dac__dac b0 b1 b2 b3 b4 vout
** GLOBAL gnd
Rresnwell@0 net@13 gnd 10k
Xr_divide@4 net@2 b2 net@1 lab_1_dac__r_divider
Xr_divide@5 net@1 b3 net@0 lab_1_dac__r_divider
Xr_divide@6 net@13 b0 net@3 lab_1_dac__r_divider
Xr_divide@7 net@0 b4 vout lab_1_dac__r_divider
Xr_divide@8 net@3 b1 net@2 lab_1_dac__r_divider
.ENDS lab_1_dac__dac

*** SUBCIRCUIT lab_1_dac__dac_gnd FROM CELL dac_gnd{sch}
.SUBCKT lab_1_dac__dac_gnd vin vout
** GLOBAL gnd
Xdac@0 gnd gnd gnd gnd vin vout lab_1_dac__dac
.ENDS lab_1_dac__dac_gnd

*** SUBCIRCUIT lab_1_dac__dac_load FROM CELL dac_load{sch}
.SUBCKT lab_1_dac__dac_load vin vout
** GLOBAL gnd
Ccap@0 gnd vout 10p
Rresnwell@0 vout gnd 10k
Xdac_gnd@1 vin vout lab_1_dac__dac_gnd
.ENDS lab_1_dac__dac_load

.global gnd

*** TOP LEVEL CELL: dac_load_sim{sch}
Xdac_cap@0 vin vout lab_1_dac__dac_load

* Spice Code nodes in cell cell 'dac_load_sim{sch}'
vin vin 0 pulse(0 2 1u 1f 1f 3u 6u)
.tran 0 2.4u 0 100p
.END
